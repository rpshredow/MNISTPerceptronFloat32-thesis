module sigmoid(
	input signed [31:0]in,
	output signed [15:0]out
);

	always @ (in) begin
		if(in >= 83886080)
			out <= 16'd4096;
		else if(in >= 83718307 && in < 83886080)
			out <= 16'd4068;
		else if(in >= 82040586 && in < 82208358)
			out <= 16'd4065;
		else if(in >= 80362864 && in < 80530636)
			out <= 16'd4062;
		else if(in >= 78685143 && in < 78852915)
			out <= 16'd4059;
		else if(in >= 77007421 && in < 77175193)
			out <= 16'd4055;
		else if(in >= 75329699 && in < 75497472)
			out <= 16'd4050;
		else if(in >= 73651978 && in < 73819750)
			out <= 16'd4046;
		else if(in >= 71974256 && in < 72142028)
			out <= 16'd4041;
		else if(in >= 70296535 && in < 70464307)
			out <= 16'd4035;
		else if(in >= 68618813 && in < 68786585)
			out <= 16'd4029;
		else if(in >= 66941091 && in < 67108864)
			out <= 16'd4022;
		else if(in >= 65263370 && in < 65431142)
			out <= 16'd4014;
		else if(in >= 63585648 && in < 63753420)
			out <= 16'd4006;
		else if(in >= 61907927 && in < 62075699)
			out <= 16'd3997;
		else if(in >= 60230205 && in < 60397977)
			out <= 16'd3987;
		else if(in >= 58552483 && in < 58720256)
			out <= 16'd3975;
		else if(in >= 56874762 && in < 57042534)
			out <= 16'd3963;
		else if(in >= 55197040 && in < 55364812)
			out <= 16'd3950;
		else if(in >= 53519319 && in < 53687091)
			out <= 16'd3935;
		else if(in >= 51841597 && in < 52009369)
			out <= 16'd3919;
		else if(in >= 50163875 && in < 50331648)
			out <= 16'd3901;
		else if(in >= 48486154 && in < 48653926)
			out <= 16'd3882;
		else if(in >= 46808432 && in < 46976204)
			out <= 16'd3861;
		else if(in >= 45130711 && in < 45298483)
			out <= 16'd3838;
		else if(in >= 43452989 && in < 43620761)
			out <= 16'd3812;
		else if(in >= 41775267 && in < 41943040)
			out <= 16'd3785;
		else if(in >= 40097546 && in < 40265318)
			out <= 16'd3755;
		else if(in >= 38419824 && in < 38587596)
			out <= 16'd3722;
		else if(in >= 36742103 && in < 36909875)
			out <= 16'd3687;
		else if(in >= 35064381 && in < 35232153)
			out <= 16'd3649;
		else if(in >= 33386659 && in < 33554432)
			out <= 16'd3607;
		else if(in >= 31708938 && in < 31876710)
			out <= 16'd3563;
		else if(in >= 30031216 && in < 30198988)
			out <= 16'd3514;
		else if(in >= 28353495 && in < 28521267)
			out <= 16'd3463;
		else if(in >= 26675773 && in < 26843545)
			out <= 16'd3407;
		else if(in >= 24998051 && in < 25165824)
			out <= 16'd3348;
		else if(in >= 23320330 && in < 23488102)
			out <= 16'd3285;
		else if(in >= 21642608 && in < 21810380)
			out <= 16'd3218;
		else if(in >= 19964887 && in < 20132659)
			out <= 16'd3147;
		else if(in >= 18287165 && in < 18454937)
			out <= 16'd3073;
		else if(in >= 16609443 && in < 16777216)
			out <= 16'd2994;
		else if(in >= 14931722 && in < 15099494)
			out <= 16'd2912;
		else if(in >= 13254000 && in < 13421772)
			out <= 16'd2826;
		else if(in >= 11576279 && in < 11744051)
			out <= 16'd2736;
		else if(in >= 9898557 && in < 10066329)
			out <= 16'd2644;
		else if(in >= 8220835 && in < 8388608)
			out <= 16'd2549;
		else if(in >= 6543114 && in < 6710886)
			out <= 16'd2452;
		else if(in >= 4865392 && in < 5033164)
			out <= 16'd2352;
		else if(in >= 3187671 && in < 3355443)
			out <= 16'd2252;
		else if(in >= 1509949 && in < 1677721)
			out <= 16'd2150;
		else if(in > -167772 && in <= 0)
			out <= 16'd2048;
		else if(in > -1845493 && in <= -1677721)
			out <= 16'd1945;
		else if(in > -3523215 && in <= -3355443)
			out <= 16'd1843;
		else if(in > -5200936 && in <= -5033164)
			out <= 16'd1743;
		else if(in > -6878658 && in <= -6710886)
			out <= 16'd1643;
		else if(in > -8556380 && in <= -8388608)
			out <= 16'd1546;
		else if(in > -10234101 && in <= -10066329)
			out <= 16'd1451;
		else if(in > -11911823 && in <= -11744051)
			out <= 16'd1359;
		else if(in > -13589544 && in <= -13421772)
			out <= 16'd1269;
		else if(in > -15267266 && in <= -15099494)
			out <= 16'd1183;
		else if(in > -16944988 && in <= -16777216)
			out <= 16'd1101;
		else if(in > -18622709 && in <= -18454937)
			out <= 16'd1022;
		else if(in > -20300431 && in <= -20132659)
			out <= 16'd948;
		else if(in > -21978152 && in <= -21810380)
			out <= 16'd877;
		else if(in > -23655874 && in <= -23488102)
			out <= 16'd810;
		else if(in > -25333596 && in <= -25165824)
			out <= 16'd747;
		else if(in > -27011317 && in <= -26843545)
			out <= 16'd688;
		else if(in > -28689039 && in <= -28521267)
			out <= 16'd632;
		else if(in > -30366760 && in <= -30198988)
			out <= 16'd581;
		else if(in > -32044482 && in <= -31876710)
			out <= 16'd532;
		else if(in > -33722204 && in <= -33554432)
			out <= 16'd488;
		else if(in > -35399925 && in <= -35232153)
			out <= 16'd446;
		else if(in > -37077647 && in <= -36909875)
			out <= 16'd408;
		else if(in > -38755368 && in <= -38587596)
			out <= 16'd373;
		else if(in > -40433090 && in <= -40265318)
			out <= 16'd340;
		else if(in > -42110812 && in <= -41943040)
			out <= 16'd310;
		else if(in > -43788533 && in <= -43620761)
			out <= 16'd283;
		else if(in > -45466255 && in <= -45298483)
			out <= 16'd257;
		else if(in > -47143976 && in <= -46976204)
			out <= 16'd234;
		else if(in > -48821698 && in <= -48653926)
			out <= 16'd213;
		else if(in > -50499420 && in <= -50331648)
			out <= 16'd194;
		else if(in > -52177141 && in <= -52009369)
			out <= 16'd176;
		else if(in > -53854863 && in <= -53687091)
			out <= 16'd160;
		else if(in > -55532584 && in <= -55364812)
			out <= 16'd145;
		else if(in > -57210306 && in <= -57042534)
			out <= 16'd132;
		else if(in > -58888028 && in <= -58720256)
			out <= 16'd120;
		else if(in > -60565749 && in <= -60397977)
			out <= 16'd108;
		else if(in > -62243471 && in <= -62075699)
			out <= 16'd98;
		else if(in > -63921192 && in <= -63753420)
			out <= 16'd89;
		else if(in > -65598914 && in <= -65431142)
			out <= 16'd81;
		else if(in > -67276636 && in <= -67108864)
			out <= 16'd73;
		else if(in > -68954357 && in <= -68786585)
			out <= 16'd66;
		else if(in > -70632079 && in <= -70464307)
			out <= 16'd60;
		else if(in > -72309800 && in <= -72142028)
			out <= 16'd54;
		else if(in > -73987522 && in <= -73819750)
			out <= 16'd49;
		else if(in > -75665244 && in <= -75497472)
			out <= 16'd45;
		else if(in > -77342965 && in <= -77175193)
			out <= 16'd40;
		else if(in > -79020687 && in <= -78852915)
			out <= 16'd36;
		else if(in > -80698408 && in <= -80530636)
			out <= 16'd33;
		else if(in > -82376130 && in <= -82208358)
			out <= 16'd30;
		else
			out <= 16'd0;
	end
endmodule
